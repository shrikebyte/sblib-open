--##############################################################################
--# File : axis_resize.vhd
--# Auth : David Gussler
--# Lang : VHDL'19
--# ============================================================================
--! AXI-Stream resizer.
--! Like most other axi stream IP, this only works properly if tkeep is
--! high on all beats except for tlast, and on tlast, upper tkeep bits should
--! be zero and lower bits should be 1.
--! When upsizing, data width, keep width, and user width should all be
--! powers of 2. Otherwise, multiplies will be inferred, greatly increasing
--! logic utilization.
--! This has a comb tready path. Insert an axi stream pipeline stage before
--! the input of this module, if needed to improve timing.
--! TODO: Change upsizer so that it will pack sparse tkeep inputs.
--##############################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.util_pkg.all;
use work.axis_pkg.all;

entity axis_resize is
  port (
    clk    : in    std_ulogic;
    srst   : in    std_ulogic;
    --
    s_axis : view s_axis_v;
    --
    m_axis : view m_axis_v;
  );
end entity;

architecture rtl of axis_resize is

  constant S_DW  : integer := s_axis.tdata'length;
  constant S_KW  : integer := s_axis.tkeep'length;
  constant S_UW  : integer := s_axis.tuser'length;
  constant S_DBW : integer := S_DW / S_KW;
  constant S_UBW : integer := S_UW / S_KW;
  constant M_DW  : integer := m_axis.tdata'length;
  constant M_KW  : integer := m_axis.tkeep'length;
  constant M_UW  : integer := m_axis.tuser'length;
  constant M_DBW : integer := M_DW / M_KW;
  constant M_UBW : integer := M_UW / M_KW;

begin

  -- ---------------------------------------------------------------------------
  assert S_DBW = M_DBW
    report "axis_resize: Input and output data byte widths must be " &
      "equal. They are implicitly defined as the ratio of data width to keep " &
      "width."
    severity error;

  assert S_UBW = M_UBW
  report "axis_resize: Input and output user byte widths must be " &
    "equal. They are implicitly defined as the ratio of user width to keep " &
    "width."
    severity error;

  prc_assert : process (clk) begin
    if rising_edge(clk) then
      assert not (s_axis.tvalid = '1' and s_axis.tlast = '1' and
        (nor s_axis.tkeep) = '1')
        report "axis_resize: Null tlast beat detected on input. At " &
          "least one tkeep bit must be set on tlast."
        severity error;

      assert not (s_axis.tvalid = '1' and not is_contig(s_axis.tkeep))
        report "axis_resize: Non-contiguous tkeep detected on input. tkeep " &
          "must be contiguous (e.g., 0001, 0011, 0111, but not 0101 or 0100)."
        severity error;
    end if;
  end process;

  -- ---------------------------------------------------------------------------
  -- Passthrough mode
  gen_resize_mode : if S_DW = M_DW generate
  begin

    s_axis.tready <= m_axis.tready;
    m_axis.tvalid <= s_axis.tvalid;
    m_axis.tlast  <= s_axis.tlast;
    m_axis.tdata  <= s_axis.tdata;
    m_axis.tkeep  <= s_axis.tkeep;
    m_axis.tuser  <= s_axis.tuser;


  -- ---------------------------------------------------------------------------
  -- Downsize mode
  elsif S_DW > M_DW generate
    constant RATIO : integer := S_DW / M_DW;
    signal last_reg  : std_ulogic_vector(RATIO - 1 downto 0);
    signal data_reg : std_ulogic_vector(S_DW-1 downto 0);
    signal user_reg : std_ulogic_vector(S_UW-1 downto 0);
    signal keep_reg : std_ulogic_vector(S_KW-1 downto 0);
    signal last_reg_shft : std_ulogic_vector(RATIO - 1 downto 0);
    signal data_reg_shft : std_ulogic_vector(S_DW-1 downto 0);
    signal user_reg_shft : std_ulogic_vector(S_UW-1 downto 0);
    signal keep_reg_shft : std_ulogic_vector(S_KW-1 downto 0);
    signal keep_reg_shft_is_zero : std_logic;
    signal tkeep_contracted : std_ulogic_vector(RATIO - 1 downto 0);

    function find_last_idx (
      vec : std_ulogic_vector
    ) return natural is
      variable tmp : natural := 0;
    begin
      for i in vec'low to vec'high loop
        if vec(i) then
          tmp := i;
        end if;
      end loop;
      return tmp;
    end function;

  begin

    -- Input is ready whenever there is room in the output buffer AND the
    -- shift register is empty.
    s_axis.tready <= (m_axis.tready or not m_axis.tvalid) and keep_reg_shft_is_zero;

    data_reg_shft <= std_ulogic_vector(shift_right(u_unsigned(data_reg), M_DW));
    user_reg_shft <= std_ulogic_vector(shift_right(u_unsigned(user_reg), M_UW));
    keep_reg_shft <= std_ulogic_vector(shift_right(u_unsigned(keep_reg), M_KW));
    last_reg_shft <= std_ulogic_vector(shift_right(u_unsigned(last_reg), 1));
    keep_reg_shft_is_zero <= and (not keep_reg_shft);

    tkeep_contracted <= contract_bits(s_axis.tkeep, M_KW);

    prc_downsize : process (clk) begin
      if rising_edge(clk) then

        if s_axis.tvalid and s_axis.tready then
          -- New wide beat at input... send the first narrow output beat.

          m_axis.tvalid <= '1';
          data_reg <= s_axis.tdata;
          user_reg <= s_axis.tuser;
          keep_reg <= s_axis.tkeep;
          last_reg <= (others=>'0');
          last_reg(find_last_idx(tkeep_contracted)) <= s_axis.tlast;

        elsif m_axis.tvalid and m_axis.tready then
          -- Shift out the narrow output data from the rest of the
          -- wide input data until the shift register is empty.

          data_reg <= data_reg_shft;
          user_reg <= user_reg_shft;
          keep_reg <= keep_reg_shft;
          last_reg <= last_reg_shft;

          if keep_reg_shft_is_zero then
            m_axis.tvalid <= '0';
          end if;

        end if;

        if srst then
          m_axis.tvalid <= '0';
          keep_reg <= (others => '0');
        end if;
      end if;
    end process;

    m_axis.tdata <= data_reg(m_axis.tdata'range);
    m_axis.tuser <= user_reg(m_axis.tuser'range);
    m_axis.tkeep <= keep_reg(m_axis.tkeep'range);
    m_axis.tlast <= last_reg(0);


  -- ---------------------------------------------------------------------------
  -- Upsize mode
  else generate
    constant CNT_MAX : integer := (M_DW / S_DW) - 1;
    signal cnt : integer range 0 to CNT_MAX;
  begin

    s_axis.tready <= m_axis.tready or not m_axis.tvalid;

    prc_upsize : process (clk) begin
      if rising_edge(clk) then
        if s_axis.tvalid and s_axis.tready then
          -- New narrow input beat

          if cnt = 0 then
            -- First narrow input beat of wide output beat
            m_axis.tkeep <= (others=>'0');
          end if;
          m_axis.tkeep(cnt * S_KW + S_KW - 1 downto cnt * S_KW) <= s_axis.tkeep;
          m_axis.tdata(cnt * S_DW + S_DW - 1 downto cnt * S_DW) <= s_axis.tdata;
          m_axis.tuser(cnt * S_UW + S_UW - 1 downto cnt * S_UW) <= s_axis.tuser;
          m_axis.tlast <= s_axis.tlast;

          if cnt = CNT_MAX or s_axis.tlast = '1' then
            m_axis.tvalid <= '1';
            cnt <= 0;
          else
            m_axis.tvalid <= '0';
            cnt <= cnt + 1;
          end if;

        elsif m_axis.tready then
          m_axis.tvalid <= '0';
        end if;

        if srst then
          m_axis.tvalid <= '0';
          cnt <= 0;
        end if;
      end if;
    end process;

  end generate;

end architecture;
